LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE MURATOV_MIPS IS

	TYPE mem_array IS ARRAY (0 TO 31) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

END MURATOV_MIPS;

PACKAGE BODY MURATOV_MIPS IS

END PACKAGE BODY;